`timescale 1ns/1ps

module 2X1tb