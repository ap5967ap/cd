module hello(A,B);

    input A;
    output B;

    not notA(B,A);


endmodule